
.include libs/LM2731Y_TRANS.LIB
.include libs/MBR0520LT1.LIB

* 1 0 3 9 9 LM2731YMF
* .SUBCKT LM2731Y_TRANS VIN SHDN_N SW FB GND
.subckt LM2731YMF 1 2 3 4 5
  XU1 5 4 1 3 2 LM2731Y_TRANS
.ends LM2731YMF

.subckt MBR0520LT 1 2
*  Dmbr0520lt1 1 2
  D1 2 1 Dmbr0520lt1
.ends MBR0520LT
