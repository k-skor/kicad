.title KiCad schematic
.include "power.cir"
.include "spice\BC548C.lib"
.include "spice\LM317A_TRANS.LIB"
XU1 VCC /TRANSISTOR_UCE /OUTPUT_14V4_P LM317A_TRANS
R1 /OUTPUT_14V4_P /TRANSISTOR_UCE 240
R2 /TRANSISTOR_UCE /OUTPUT_14V4_N 2.55k
R3 /OUTPUT_14V4_N 0 1
Q1 /TRANSISTOR_UCE /OUTPUT_14V4_N 0 BC548C
XP1 VCC 0 PWR_IN
R4 /OUTPUT_14V4_P /OUTPUT_14V4_N 30
C1 VCC 0 0.1u
C2 /OUTPUT_14V4_P /OUTPUT_14V4_N 1u
.tran 10us 1ms uic 
.end
