* /home/krzy0s/snap/kicad-snap/common/opamp/opamp2.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: nie, 19 lis 2017, 22:18:32

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

.include components.cir

* Sheet Name: /
XU1  ? 8 4 3 ? 6 1 LM741		
R1  8 0 1K		
R2  6 8 2K		
XP1  1 0 3 PWR_IN		
XJ1  4 0 SRC_IN		

.op

.end
