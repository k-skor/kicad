.subckt PWR_IN 1 2
  Vin 1 2 18
.ends PWR_IN
