.title KiCad schematic
.include common.cir
.include "libs/LM2731Y_TRANS.LIB"
.include "libs/MBR0520LT1.LIB"
*.include "power.cir"
C1 VCC 0 2u2
C2 /INPUT_18V Net-_C2-Pad2_ 150p
C3 /INPUT_18V 0 4u7
R1 Net-_C2-Pad2_ 0 13k3
R2 /INPUT_18V Net-_C2-Pad2_ 181k3
R3 0 /INPUT_18V 180
XU1 Net-_D1-Pad2_ 0 Net-_C2-Pad2_ VCC VCC LM2731Y_TRANS
D1 Net-_D1-Pad2_ /INPUT_18V Dmbr0520lt1
*XP1 VCC 0 PWR_IN
L1 VCC Net-_D1-Pad2_ 10u
Vcc VCC 0 12
.tran 10us 500us uic
.end
