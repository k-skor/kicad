.title KiCad schematic
.include "libs/BC548C.lib"
.include "libs/LM317A_TRANS.LIB"
.include "power.cir"
XU1 VCC Net-_Q1-Pad1_ /OUTPUT_14V4_P LM317A_TRANS
R1 /OUTPUT_14V4_P Net-_Q1-Pad1_ 240
R2 Net-_Q1-Pad1_ /OUTPUT_14V4_N 3k117
R3 /OUTPUT_14V4_N 0 1
Q1 Net-_Q1-Pad1_ /OUTPUT_14V4_N 0 BC548C
XP1 VCC 0 PWR_IN
R4 /OUTPUT_14V4_P /OUTPUT_14V4_N 30
.tran 10us 1ms uic
.end
