.subckt PWR_IN 1 2
  Vin 1 2 12
.ends PWR_IN
